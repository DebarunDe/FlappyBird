module Bird (

);



endmodule
