module FlappyBird (


);



endmodule 